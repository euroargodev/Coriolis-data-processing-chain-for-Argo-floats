netcdf ArgoV2MergedProf_V1.0 {
dimensions:
	DATE_TIME = 14 ;
	STRING256 = 256 ;
	STRING64 = 64 ;
	STRING32 = 32 ;
	STRING8 = 8 ;
	STRING4 = 4 ;
	STRING2 = 2 ;
	N_PROF = 1 ;
	N_PARAM = 1 ;
	N_LEVELS = 1 ;
	N_CALIB = 1 ;
variables:
	char DATA_TYPE(STRING32) ;
		DATA_TYPE:long_name = "Data type" ;
		DATA_TYPE:conventions = "Argo reference table 1" ;
		DATA_TYPE:_FillValue = " " ;
	char FORMAT_VERSION(STRING4) ;
		FORMAT_VERSION:long_name = "File format version" ;
		FORMAT_VERSION:_FillValue = " " ;
	char HANDBOOK_VERSION(STRING4) ;
		HANDBOOK_VERSION:long_name = "Data handbook version" ;
		HANDBOOK_VERSION:_FillValue = " " ;
	char REFERENCE_DATE_TIME(DATE_TIME) ;
		REFERENCE_DATE_TIME:long_name = "Date of reference for Julian days" ;
		REFERENCE_DATE_TIME:conventions = "YYYYMMDDHHMISS" ;
		REFERENCE_DATE_TIME:_FillValue = " " ;
	char DATE_CREATION(DATE_TIME) ;
		DATE_CREATION:long_name = "Date of file creation" ;
		DATE_CREATION:conventions = "YYYYMMDDHHMISS" ;
		DATE_CREATION:_FillValue = " " ;
	char DATE_UPDATE(DATE_TIME) ;
		DATE_UPDATE:long_name = "Date of update of this file" ;
		DATE_UPDATE:conventions = "YYYYMMDDHHMISS" ;
		DATE_UPDATE:_FillValue = " " ;
	char PLATFORM_NUMBER(N_PROF, STRING8) ;
		PLATFORM_NUMBER:long_name = "Float unique identifier" ;
		PLATFORM_NUMBER:conventions = "WMO float identifier : A9IIIII" ;
		PLATFORM_NUMBER:_FillValue = " " ;
	char PROJECT_NAME(N_PROF, STRING64) ;
		PROJECT_NAME:long_name = "Name of the project" ;
		PROJECT_NAME:_FillValue = " " ;
	char PI_NAME(N_PROF, STRING64) ;
		PI_NAME:long_name = "Name of the principal investigator" ;
		PI_NAME:_FillValue = " " ;
	char STATION_PARAMETERS(N_PROF, N_PARAM, STRING64) ;
		STATION_PARAMETERS:long_name = "List of available parameters for the station" ;
		STATION_PARAMETERS:conventions = "Argo reference table 3" ;
		STATION_PARAMETERS:_FillValue = " " ;
	int CYCLE_NUMBER(N_PROF) ;
		CYCLE_NUMBER:long_name = "Float cycle number" ;
		CYCLE_NUMBER:conventions = "0...N, 0 : launch cycle (if exists), 1 : first complete cycle" ;
		CYCLE_NUMBER:_FillValue = 99999 ;
	char DIRECTION(N_PROF) ;
		DIRECTION:long_name = "Direction of the station profiles" ;
		DIRECTION:conventions = "A: ascending profiles, D: descending profiles" ;
		DIRECTION:_FillValue = " " ;
	char DATA_CENTRE(N_PROF, STRING2) ;
		DATA_CENTRE:long_name = "Data centre in charge of float data processing" ;
		DATA_CENTRE:conventions = "Argo reference table 4" ;
		DATA_CENTRE:_FillValue = " " ;
	char PARAMETER_DATA_MODE(N_PROF, N_PARAM) ;
		PARAMETER_DATA_MODE:long_name = "Delayed mode or real time data" ;
		PARAMETER_DATA_MODE:conventions = "R : real time; D : delayed mode; A : real time with adjustment" ;
		PARAMETER_DATA_MODE:_FillValue = " " ;
	char PLATFORM_TYPE(N_PROF, STRING32) ;
		PLATFORM_TYPE:long_name = "Type of float" ;
		PLATFORM_TYPE:conventions = "Argo reference table 23" ;
		PLATFORM_TYPE:_FillValue = " " ;
	char FLOAT_SERIAL_NO(N_PROF, STRING32) ;
		FLOAT_SERIAL_NO:long_name = "Serial number of the float" ;
		FLOAT_SERIAL_NO:_FillValue = " " ;
	char FIRMWARE_VERSION(N_PROF, STRING32) ;
		FIRMWARE_VERSION:long_name = "Instrument firmware version" ;
		FIRMWARE_VERSION:_FillValue = " " ;
	char WMO_INST_TYPE(N_PROF, STRING4) ;
		WMO_INST_TYPE:long_name = "Coded instrument type" ;
		WMO_INST_TYPE:conventions = "Argo reference table 8" ;
		WMO_INST_TYPE:_FillValue = " " ;
	double JULD(N_PROF) ;
		JULD:long_name = "Julian day (UTC) of the station relative to REFERENCE_DATE_TIME" ;
		JULD:standard_name = "time" ;
		JULD:units = "days since 1950-01-01 00:00:00 UTC" ;
		JULD:conventions = "Relative julian days with decimal part (as parts of day)" ;
		JULD:_FillValue = 999999. ;
		JULD:axis = "T" ;
	char JULD_QC(N_PROF) ;
		JULD_QC:long_name = "Quality on date and time" ;
		JULD_QC:conventions = "Argo reference table 2" ;
		JULD_QC:_FillValue = " " ;
	double JULD_LOCATION(N_PROF) ;
		JULD_LOCATION:long_name = "Julian day (UTC) of the location relative to REFERENCE_DATE_TIME" ;
		JULD_LOCATION:units = "days since 1950-01-01 00:00:00 UTC" ;
		JULD_LOCATION:conventions = "Relative julian days with decimal part (as parts of day)" ;
		JULD_LOCATION:_FillValue = 999999. ;
	double LATITUDE(N_PROF) ;
		LATITUDE:long_name = "Latitude of the station, best estimate" ;
		LATITUDE:standard_name = "latitude" ;
		LATITUDE:units = "degree_north" ;
		LATITUDE:_FillValue = 99999. ;
		LATITUDE:valid_min = -90. ;
		LATITUDE:valid_max = 90. ;
		LATITUDE:axis = "Y" ;
	double LONGITUDE(N_PROF) ;
		LONGITUDE:long_name = "Longitude of the station, best estimate" ;
		LONGITUDE:standard_name = "longitude" ;
		LONGITUDE:units = "degree_east" ;
		LONGITUDE:_FillValue = 99999. ;
		LONGITUDE:valid_min = -180. ;
		LONGITUDE:valid_max = 180. ;
		LONGITUDE:axis = "X" ;
	char POSITION_QC(N_PROF) ;
		POSITION_QC:long_name = "Quality on position (latitude and longitude)" ;
		POSITION_QC:conventions = "Argo reference table 2" ;
		POSITION_QC:_FillValue = " " ;
	char POSITIONING_SYSTEM(N_PROF, STRING8) ;
		POSITIONING_SYSTEM:long_name = "Positioning system" ;
		POSITIONING_SYSTEM:_FillValue = " " ;
	int CONFIG_MISSION_NUMBER(N_PROF) ;
		CONFIG_MISSION_NUMBER:long_name = "Unique number denoting the missions performed by the float" ;
		CONFIG_MISSION_NUMBER:conventions = "1...N, 1 : first complete mission" ;
		CONFIG_MISSION_NUMBER:_FillValue = 99999 ;
	char PARAMETER(N_PROF, N_CALIB, N_PARAM, STRING64) ;
		PARAMETER:long_name = "List of parameters with calibration information" ;
		PARAMETER:conventions = "Argo reference table 3" ;
		PARAMETER:_FillValue = " " ;
	char SCIENTIFIC_CALIB_EQUATION(N_PROF, N_CALIB, N_PARAM, STRING256) ;
		SCIENTIFIC_CALIB_EQUATION:long_name = "Calibration equation for this parameter" ;
		SCIENTIFIC_CALIB_EQUATION:_FillValue = " " ;
	char SCIENTIFIC_CALIB_COEFFICIENT(N_PROF, N_CALIB, N_PARAM, STRING256) ;
		SCIENTIFIC_CALIB_COEFFICIENT:long_name = "Calibration coefficients for this equation" ;
		SCIENTIFIC_CALIB_COEFFICIENT:_FillValue = " " ;
	char SCIENTIFIC_CALIB_COMMENT(N_PROF, N_CALIB, N_PARAM, STRING256) ;
		SCIENTIFIC_CALIB_COMMENT:long_name = "Comment applying to this parameter calibration" ;
		SCIENTIFIC_CALIB_COMMENT:_FillValue = " " ;
	char SCIENTIFIC_CALIB_DATE(N_PROF, N_CALIB, N_PARAM, DATE_TIME) ;
		SCIENTIFIC_CALIB_DATE:long_name = "Date of calibration" ;
		SCIENTIFIC_CALIB_DATE:conventions = "YYYYMMDDHHMISS" ;
		SCIENTIFIC_CALIB_DATE:_FillValue = " " ;
		
// global attributes:
		:title = "" ;
		:institution = "" ;
		:source = "" ;
		:history = "" ;
		:references = "" ;
		:user_manual_version = "" ;
		:Conventions = "" ;
		:featureType = "" ;
data:

 DATA_TYPE = " " ;

 FORMAT_VERSION = " " ;

 HANDBOOK_VERSION = " " ;

 REFERENCE_DATE_TIME = " " ;

 DATE_CREATION = " " ;

 DATE_UPDATE = " " ;

 PLATFORM_NUMBER = " " ;

 PROJECT_NAME = " " ;

 PI_NAME = " " ;

 STATION_PARAMETERS = " " ;

 CYCLE_NUMBER = _ ;

 DIRECTION = " " ;

 DATA_CENTRE = " " ;

 PARAMETER_DATA_MODE = " " ;

 PLATFORM_TYPE = " " ;

 FLOAT_SERIAL_NO = " " ;

 FIRMWARE_VERSION = " " ;

 WMO_INST_TYPE = " " ;

 JULD = _ ;

 JULD_QC = " " ;

 JULD_LOCATION = _ ;

 LATITUDE = _ ;

 LONGITUDE = _ ;

 POSITION_QC = " " ;

 POSITIONING_SYSTEM = " " ;

 CONFIG_MISSION_NUMBER = _ ;

 PARAMETER = "" ;

 SCIENTIFIC_CALIB_EQUATION = "" ;

 SCIENTIFIC_CALIB_COMMENT = "" ;

 SCIENTIFIC_CALIB_DATE = "" ;
}
