version https://git-lfs.github.com/spec/v1
oid sha256:02b490a1d61d3a677dcd7002e617e6ba91448bc0c91742ff17b9e10ade3b2bef
size 7554
