version https://git-lfs.github.com/spec/v1
oid sha256:d84628fa88e577b6a901abb073f40bfb243cd27818fd85c0f7ff0f5dc96d48a4
size 7547
